`timescale 1ns / 1ps

module and2(output y_out, input a, b);
    and (y_out, a, b);
endmodule